VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_urish_skullfet
  CLASS BLOCK ;
  FOREIGN tt_um_urish_skullfet ;
  ORIGIN 0.000 0.000 ;
  SIZE 157.320 BY 111.520 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 12.315 2.480 13.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 22.315 2.480 23.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 32.315 2.480 33.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 42.315 2.480 43.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 52.315 2.480 53.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 62.315 2.480 63.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 72.315 2.480 73.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.315 2.480 83.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 92.315 2.480 93.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 102.315 2.480 103.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 112.315 2.480 113.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 122.315 2.480 123.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 132.315 2.480 133.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 142.315 2.480 143.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 152.315 2.480 153.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.260 24.240 5.860 68.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 7.315 2.480 8.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 17.315 2.480 18.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.315 2.480 28.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 37.315 2.480 38.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.315 2.480 48.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.315 2.480 58.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 67.315 2.480 68.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 77.315 2.480 78.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 87.315 2.480 88.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.315 2.480 98.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 107.315 2.480 108.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 117.315 2.480 118.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 127.315 2.480 128.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 137.315 2.480 138.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 147.315 2.480 148.915 109.040 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.630 110.520 134.930 111.520 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 131.870 110.520 132.170 111.520 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 129.110 110.520 129.410 111.520 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 126.350 110.520 126.650 111.520 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 123.590 110.520 123.890 111.520 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 120.830 110.520 121.130 111.520 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 110.520 118.370 111.520 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 115.310 110.520 115.610 111.520 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.550 110.520 112.850 111.520 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 109.790 110.520 110.090 111.520 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 110.520 107.330 111.520 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 104.270 110.520 104.570 111.520 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 101.510 110.520 101.810 111.520 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 98.750 110.520 99.050 111.520 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 110.520 96.290 111.520 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.230 110.520 93.530 111.520 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.470 110.520 90.770 111.520 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 87.710 110.520 88.010 111.520 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 40.790 110.520 41.090 111.520 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 38.030 110.520 38.330 111.520 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 35.270 110.520 35.570 111.520 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 32.510 110.520 32.810 111.520 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 29.750 110.520 30.050 111.520 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 26.990 110.520 27.290 111.520 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 24.230 110.520 24.530 111.520 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 62.870 110.520 63.170 111.520 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 60.110 110.520 60.410 111.520 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 57.350 110.520 57.650 111.520 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 54.590 110.520 54.890 111.520 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 51.830 110.520 52.130 111.520 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 49.070 110.520 49.370 111.520 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 46.310 110.520 46.610 111.520 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 43.550 110.520 43.850 111.520 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 84.950 110.520 85.250 111.520 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 82.190 110.520 82.490 111.520 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 79.430 110.520 79.730 111.520 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 76.670 110.520 76.970 111.520 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 73.910 110.520 74.210 111.520 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 71.150 110.520 71.450 111.520 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 68.390 110.520 68.690 111.520 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 65.630 110.520 65.930 111.520 ;
    END
  END uo_out[7]
  OBS
      LAYER nwell ;
        RECT 2.570 107.385 154.750 108.990 ;
        RECT 2.570 101.945 154.750 104.775 ;
        RECT 2.570 96.505 154.750 99.335 ;
        RECT 2.570 91.065 154.750 93.895 ;
        RECT 2.570 85.625 154.750 88.455 ;
        RECT 2.570 80.185 154.750 83.015 ;
        RECT 2.570 74.745 154.750 77.575 ;
        RECT 2.570 69.305 154.750 72.135 ;
        RECT 2.570 65.090 154.750 66.695 ;
        RECT 2.570 63.865 20.430 65.090 ;
        RECT 2.570 58.425 20.430 61.255 ;
        RECT 2.570 52.985 20.430 55.815 ;
        RECT 2.570 49.150 20.430 50.375 ;
        RECT 2.570 47.545 154.750 49.150 ;
        RECT 2.570 42.105 20.430 44.935 ;
        RECT 2.570 36.665 20.430 39.495 ;
        RECT 2.570 31.225 20.430 34.055 ;
        RECT 2.570 27.390 20.430 28.615 ;
        RECT 2.570 25.785 154.750 27.390 ;
        RECT 2.570 20.345 154.750 23.175 ;
        RECT 2.570 14.905 154.750 17.735 ;
        RECT 2.570 9.465 154.750 12.295 ;
        RECT 2.570 4.025 154.750 6.855 ;
      LAYER li1 ;
        RECT 2.760 2.635 154.560 108.885 ;
      LAYER met1 ;
        RECT 2.760 2.480 154.560 109.040 ;
      LAYER met2 ;
        RECT 4.290 2.535 153.885 110.005 ;
      LAYER met3 ;
        RECT 4.270 2.555 153.905 109.985 ;
      LAYER met4 ;
        RECT 22.170 110.120 23.830 110.520 ;
        RECT 24.930 110.120 26.590 110.520 ;
        RECT 27.690 110.120 29.350 110.520 ;
        RECT 30.450 110.120 32.110 110.520 ;
        RECT 33.210 110.120 34.870 110.520 ;
        RECT 35.970 110.120 37.630 110.520 ;
        RECT 38.730 110.120 40.390 110.520 ;
        RECT 41.490 110.120 43.150 110.520 ;
        RECT 44.250 110.120 45.910 110.520 ;
        RECT 47.010 110.120 48.670 110.520 ;
        RECT 49.770 110.120 51.430 110.520 ;
        RECT 52.530 110.120 54.190 110.520 ;
        RECT 55.290 110.120 56.950 110.520 ;
        RECT 58.050 110.120 59.710 110.520 ;
        RECT 60.810 110.120 62.470 110.520 ;
        RECT 63.570 110.120 65.230 110.520 ;
        RECT 66.330 110.120 67.990 110.520 ;
        RECT 69.090 110.120 70.750 110.520 ;
        RECT 71.850 110.120 73.510 110.520 ;
        RECT 74.610 110.120 76.270 110.520 ;
        RECT 77.370 110.120 79.030 110.520 ;
        RECT 80.130 110.120 81.790 110.520 ;
        RECT 82.890 110.120 84.550 110.520 ;
        RECT 85.650 110.120 87.310 110.520 ;
        RECT 88.410 110.120 90.070 110.520 ;
        RECT 91.170 110.120 92.830 110.520 ;
        RECT 93.930 110.120 95.590 110.520 ;
        RECT 96.690 110.120 98.350 110.520 ;
        RECT 99.450 110.120 101.110 110.520 ;
        RECT 102.210 110.120 103.870 110.520 ;
        RECT 104.970 110.120 106.630 110.520 ;
        RECT 107.730 110.120 109.390 110.520 ;
        RECT 110.490 110.120 112.150 110.520 ;
        RECT 113.250 110.120 114.910 110.520 ;
        RECT 116.010 110.120 117.670 110.520 ;
        RECT 118.770 110.120 120.430 110.520 ;
        RECT 121.530 110.120 123.190 110.520 ;
        RECT 124.290 110.120 125.950 110.520 ;
        RECT 127.050 110.120 128.710 110.520 ;
        RECT 129.810 110.120 130.345 110.520 ;
        RECT 21.455 109.440 130.345 110.120 ;
        RECT 21.455 108.975 21.915 109.440 ;
        RECT 24.315 108.975 26.915 109.440 ;
        RECT 29.315 108.975 31.915 109.440 ;
        RECT 34.315 108.975 36.915 109.440 ;
        RECT 39.315 108.975 41.915 109.440 ;
        RECT 44.315 108.975 46.915 109.440 ;
        RECT 49.315 108.975 51.915 109.440 ;
        RECT 54.315 108.975 56.915 109.440 ;
        RECT 59.315 108.975 61.915 109.440 ;
        RECT 64.315 108.975 66.915 109.440 ;
        RECT 69.315 108.975 71.915 109.440 ;
        RECT 74.315 108.975 76.915 109.440 ;
        RECT 79.315 108.975 81.915 109.440 ;
        RECT 84.315 108.975 86.915 109.440 ;
        RECT 89.315 108.975 91.915 109.440 ;
        RECT 94.315 108.975 96.915 109.440 ;
        RECT 99.315 108.975 101.915 109.440 ;
        RECT 104.315 108.975 106.915 109.440 ;
        RECT 109.315 108.975 111.915 109.440 ;
        RECT 114.315 108.975 116.915 109.440 ;
        RECT 119.315 108.975 121.915 109.440 ;
        RECT 124.315 108.975 126.915 109.440 ;
        RECT 129.315 108.975 130.345 109.440 ;
  END
END tt_um_urish_skullfet
END LIBRARY

