VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_urish_ringosc_cnt
  CLASS BLOCK ;
  FOREIGN tt_um_urish_ringosc_cnt ;
  ORIGIN 0.000 0.000 ;
  SIZE 168.360 BY 111.520 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 109.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 109.040 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 145.670 110.520 145.970 111.520 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 148.430 110.520 148.730 111.520 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 142.910 110.520 143.210 111.520 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 140.150 110.520 140.450 111.520 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 134.630 110.520 134.930 111.520 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 131.870 110.520 132.170 111.520 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 129.110 110.520 129.410 111.520 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 126.350 110.520 126.650 111.520 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 123.590 110.520 123.890 111.520 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 120.830 110.520 121.130 111.520 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 110.520 118.370 111.520 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 115.310 110.520 115.610 111.520 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.550 110.520 112.850 111.520 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 109.790 110.520 110.090 111.520 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 110.520 107.330 111.520 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 104.270 110.520 104.570 111.520 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 101.510 110.520 101.810 111.520 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 98.750 110.520 99.050 111.520 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 51.830 110.520 52.130 111.520 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 49.070 110.520 49.370 111.520 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 46.310 110.520 46.610 111.520 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 43.550 110.520 43.850 111.520 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 40.790 110.520 41.090 111.520 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 38.030 110.520 38.330 111.520 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 35.270 110.520 35.570 111.520 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 32.510 110.520 32.810 111.520 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 73.910 110.520 74.210 111.520 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 71.150 110.520 71.450 111.520 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 68.390 110.520 68.690 111.520 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 65.630 110.520 65.930 111.520 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 62.870 110.520 63.170 111.520 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 60.110 110.520 60.410 111.520 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 57.350 110.520 57.650 111.520 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 54.590 110.520 54.890 111.520 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 95.990 110.520 96.290 111.520 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 93.230 110.520 93.530 111.520 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 90.470 110.520 90.770 111.520 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 87.710 110.520 88.010 111.520 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 84.950 110.520 85.250 111.520 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 82.190 110.520 82.490 111.520 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 79.430 110.520 79.730 111.520 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 76.670 110.520 76.970 111.520 ;
    END
  END uo_out[7]
  OBS
      LAYER nwell ;
        RECT 2.570 107.385 165.790 108.990 ;
        RECT 2.570 101.945 165.790 104.775 ;
        RECT 2.570 96.505 165.790 99.335 ;
        RECT 2.570 91.065 165.790 93.895 ;
        RECT 2.570 85.625 165.790 88.455 ;
        RECT 2.570 80.185 165.790 83.015 ;
        RECT 2.570 74.745 165.790 77.575 ;
        RECT 2.570 69.305 165.790 72.135 ;
        RECT 2.570 63.865 165.790 66.695 ;
        RECT 2.570 58.425 165.790 61.255 ;
        RECT 2.570 52.985 165.790 55.815 ;
        RECT 2.570 47.545 165.790 50.375 ;
        RECT 2.570 42.105 165.790 44.935 ;
        RECT 2.570 36.665 165.790 39.495 ;
        RECT 2.570 31.225 165.790 34.055 ;
        RECT 2.570 25.785 165.790 28.615 ;
        RECT 2.570 20.345 165.790 23.175 ;
        RECT 2.570 14.905 165.790 17.735 ;
        RECT 2.570 9.465 165.790 12.295 ;
        RECT 2.570 4.025 165.790 6.855 ;
      LAYER li1 ;
        RECT 2.760 2.635 165.600 108.885 ;
      LAYER met1 ;
        RECT 2.760 2.480 165.600 110.120 ;
      LAYER met2 ;
        RECT 5.160 2.535 160.440 110.150 ;
      LAYER met3 ;
        RECT 18.290 2.555 146.675 109.985 ;
      LAYER met4 ;
        RECT 33.210 110.120 34.870 111.170 ;
        RECT 35.970 110.120 37.630 111.170 ;
        RECT 38.730 110.120 40.390 111.170 ;
        RECT 41.490 110.120 43.150 111.170 ;
        RECT 44.250 110.120 45.910 111.170 ;
        RECT 47.010 110.120 48.670 111.170 ;
        RECT 49.770 110.120 51.430 111.170 ;
        RECT 52.530 110.120 54.190 111.170 ;
        RECT 55.290 110.120 56.950 111.170 ;
        RECT 58.050 110.120 59.710 111.170 ;
        RECT 60.810 110.120 62.470 111.170 ;
        RECT 63.570 110.120 65.230 111.170 ;
        RECT 66.330 110.120 67.990 111.170 ;
        RECT 69.090 110.120 70.750 111.170 ;
        RECT 71.850 110.120 73.510 111.170 ;
        RECT 74.610 110.120 76.270 111.170 ;
        RECT 77.370 110.120 79.030 111.170 ;
        RECT 80.130 110.120 81.790 111.170 ;
        RECT 82.890 110.120 84.550 111.170 ;
        RECT 85.650 110.120 87.310 111.170 ;
        RECT 88.410 110.120 90.070 111.170 ;
        RECT 91.170 110.120 92.830 111.170 ;
        RECT 93.930 110.120 95.590 111.170 ;
        RECT 96.690 110.120 98.350 111.170 ;
        RECT 99.450 110.120 101.110 111.170 ;
        RECT 102.210 110.120 103.870 111.170 ;
        RECT 104.970 110.120 106.630 111.170 ;
        RECT 107.730 110.120 109.390 111.170 ;
        RECT 110.490 110.120 112.150 111.170 ;
        RECT 113.250 110.120 114.910 111.170 ;
        RECT 116.010 110.120 117.670 111.170 ;
        RECT 118.770 110.120 120.430 111.170 ;
        RECT 121.530 110.120 123.190 111.170 ;
        RECT 124.290 110.120 125.950 111.170 ;
        RECT 127.050 110.120 128.710 111.170 ;
        RECT 129.810 110.120 131.470 111.170 ;
        RECT 132.570 110.120 134.230 111.170 ;
        RECT 135.330 110.120 136.990 111.170 ;
        RECT 138.090 110.120 139.750 111.170 ;
        RECT 140.850 110.120 142.305 111.170 ;
        RECT 32.495 109.440 142.305 110.120 ;
        RECT 32.495 106.255 94.680 109.440 ;
        RECT 97.080 106.255 142.305 109.440 ;
  END
END tt_um_urish_ringosc_cnt
END LIBRARY

