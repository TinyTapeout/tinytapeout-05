VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_matt_divider_test
  CLASS BLOCK ;
  FOREIGN tt_um_matt_divider_test ;
  ORIGIN 0.000 0.000 ;
  SIZE 157.320 BY 111.520 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.630 110.520 134.930 111.520 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 131.870 110.520 132.170 111.520 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 110.520 129.410 111.520 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 126.350 110.520 126.650 111.520 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 123.590 110.520 123.890 111.520 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 120.830 110.520 121.130 111.520 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 110.520 118.370 111.520 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 115.310 110.520 115.610 111.520 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.550 110.520 112.850 111.520 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 109.790 110.520 110.090 111.520 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 110.520 107.330 111.520 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 104.270 110.520 104.570 111.520 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 101.510 110.520 101.810 111.520 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 98.750 110.520 99.050 111.520 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 110.520 96.290 111.520 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.230 110.520 93.530 111.520 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.470 110.520 90.770 111.520 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 87.710 110.520 88.010 111.520 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 110.520 41.090 111.520 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.030 110.520 38.330 111.520 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.270 110.520 35.570 111.520 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 32.510 110.520 32.810 111.520 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 110.520 30.050 111.520 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.990 110.520 27.290 111.520 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.230 110.520 24.530 111.520 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 110.520 63.170 111.520 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 60.110 110.520 60.410 111.520 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 57.350 110.520 57.650 111.520 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 54.590 110.520 54.890 111.520 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 110.520 52.130 111.520 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.070 110.520 49.370 111.520 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.310 110.520 46.610 111.520 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 43.550 110.520 43.850 111.520 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 110.520 85.250 111.520 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 82.190 110.520 82.490 111.520 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 79.430 110.520 79.730 111.520 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 76.670 110.520 76.970 111.520 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 110.520 74.210 111.520 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 71.150 110.520 71.450 111.520 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.390 110.520 68.690 111.520 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 65.630 110.520 65.930 111.520 ;
    END
  END uo_out[7]
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 38.360 2.990 63.950 106.180 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 113.050 4.240 138.640 107.430 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 75.340 93.730 75.670 93.900 ;
        RECT 75.880 93.730 76.210 93.900 ;
        RECT 76.420 93.730 76.750 93.900 ;
        RECT 76.960 93.730 77.290 93.900 ;
        RECT 75.420 91.915 75.590 93.730 ;
        RECT 75.960 91.915 76.130 93.730 ;
        RECT 76.500 91.915 76.670 93.730 ;
        RECT 77.040 91.915 77.210 93.730 ;
        RECT 75.420 88.280 75.590 90.095 ;
        RECT 75.960 88.280 76.130 90.095 ;
        RECT 76.500 88.280 76.670 90.095 ;
        RECT 77.040 88.280 77.210 90.095 ;
        RECT 75.340 88.110 75.670 88.280 ;
        RECT 75.880 88.110 76.210 88.280 ;
        RECT 76.420 88.110 76.750 88.280 ;
        RECT 76.960 88.110 77.290 88.280 ;
      LAYER mcon ;
        RECT 75.420 88.110 75.590 90.095 ;
        RECT 75.960 88.110 76.130 90.095 ;
        RECT 76.500 88.110 76.670 90.095 ;
        RECT 77.040 88.110 77.210 90.095 ;
      LAYER met1 ;
        RECT 71.170 97.660 72.930 99.690 ;
        RECT 75.280 98.330 77.040 99.690 ;
        RECT 75.280 97.660 76.790 98.330 ;
        RECT 83.940 97.740 85.700 99.770 ;
        RECT 71.500 89.380 72.850 97.660 ;
        RECT 75.360 96.130 76.760 97.660 ;
        RECT 84.190 97.140 85.400 97.740 ;
        RECT 87.700 97.610 89.460 99.640 ;
        RECT 75.380 93.960 75.980 96.130 ;
        RECT 84.190 95.150 85.450 97.140 ;
        RECT 87.990 96.180 89.380 97.610 ;
        RECT 75.380 93.920 76.160 93.960 ;
        RECT 76.470 93.930 76.700 93.960 ;
        RECT 77.010 93.930 77.240 93.960 ;
        RECT 75.360 91.860 76.170 93.920 ;
        RECT 76.450 93.710 77.260 93.930 ;
        RECT 84.360 93.710 85.370 95.150 ;
        RECT 76.450 92.860 85.390 93.710 ;
        RECT 76.450 91.870 77.260 92.860 ;
        RECT 84.360 92.660 85.370 92.860 ;
        RECT 75.390 91.855 75.620 91.860 ;
        RECT 75.930 91.855 76.160 91.860 ;
        RECT 76.470 91.855 76.700 91.870 ;
        RECT 77.010 91.855 77.240 91.870 ;
        RECT 75.390 90.080 75.620 90.155 ;
        RECT 75.930 90.130 76.160 90.155 ;
        RECT 76.470 90.130 76.700 90.155 ;
        RECT 77.010 90.140 77.240 90.155 ;
        RECT 73.870 89.380 75.690 90.080 ;
        RECT 71.500 88.220 75.690 89.380 ;
        RECT 71.500 87.960 72.850 88.220 ;
        RECT 73.870 88.000 75.690 88.220 ;
        RECT 75.930 89.050 76.740 90.130 ;
        RECT 77.010 89.450 78.850 90.140 ;
        RECT 87.990 89.450 89.340 96.180 ;
        RECT 75.930 88.050 76.760 89.050 ;
        RECT 77.010 88.060 89.340 89.450 ;
        RECT 77.010 88.050 77.240 88.060 ;
        RECT 76.060 87.290 76.760 88.050 ;
        RECT 78.200 88.010 89.340 88.060 ;
        RECT 87.990 87.880 89.340 88.010 ;
        RECT 76.060 86.320 82.160 87.290 ;
        RECT 76.060 86.260 76.760 86.320 ;
      LAYER via ;
        RECT 71.320 97.940 72.780 99.320 ;
        RECT 75.480 98.080 76.740 99.370 ;
        RECT 84.140 98.260 85.400 99.550 ;
        RECT 88.000 98.160 89.260 99.450 ;
        RECT 81.170 86.470 81.940 87.140 ;
      LAYER met2 ;
        RECT 70.700 97.440 73.350 99.840 ;
        RECT 75.010 97.610 77.660 100.010 ;
        RECT 79.440 98.780 82.090 100.060 ;
        RECT 79.440 97.660 82.120 98.780 ;
        RECT 83.860 97.860 86.510 100.260 ;
        RECT 87.670 97.890 90.320 100.290 ;
        RECT 80.910 86.260 82.120 97.660 ;
      LAYER via2 ;
        RECT 71.080 97.880 72.780 99.440 ;
        RECT 75.580 98.200 77.290 99.750 ;
        RECT 79.760 98.150 81.470 99.700 ;
        RECT 84.000 98.070 85.600 99.930 ;
        RECT 88.000 98.010 89.980 99.820 ;
      LAYER met3 ;
        RECT 76.410 109.070 76.790 109.080 ;
        RECT 87.140 109.070 87.460 109.110 ;
        RECT 76.410 108.770 87.460 109.070 ;
        RECT 76.410 108.760 76.790 108.770 ;
        RECT 87.140 108.730 87.460 108.770 ;
        RECT 70.850 97.630 73.090 99.670 ;
        RECT 74.930 97.370 77.590 100.010 ;
        RECT 79.320 97.600 81.960 100.290 ;
        RECT 83.300 97.680 86.190 100.520 ;
        RECT 87.770 97.830 90.240 100.130 ;
        RECT 101.040 88.830 101.610 104.140 ;
        RECT 65.930 52.530 87.790 72.930 ;
        RECT 88.990 52.530 110.850 72.930 ;
        RECT 65.930 30.930 87.790 51.330 ;
        RECT 88.990 30.930 110.850 51.330 ;
        RECT 65.930 9.330 87.790 29.730 ;
        RECT 88.990 9.330 110.850 29.730 ;
      LAYER via3 ;
        RECT 76.440 108.760 76.760 109.080 ;
        RECT 87.140 108.760 87.460 109.080 ;
        RECT 101.200 103.810 101.520 104.130 ;
        RECT 71.070 97.850 72.690 99.340 ;
        RECT 75.500 97.860 77.260 99.750 ;
        RECT 79.710 97.940 81.470 99.830 ;
        RECT 83.480 97.910 85.990 100.390 ;
        RECT 88.000 98.010 89.980 99.820 ;
        RECT 101.205 88.895 101.525 89.215 ;
        RECT 87.370 52.670 87.690 72.790 ;
        RECT 110.430 52.670 110.750 72.790 ;
        RECT 87.370 31.070 87.690 51.190 ;
        RECT 110.430 31.070 110.750 51.190 ;
        RECT 87.370 9.470 87.690 29.590 ;
        RECT 110.430 9.470 110.750 29.590 ;
      LAYER met4 ;
        RECT 76.660 110.520 76.670 110.970 ;
        RECT 79.050 110.520 79.430 110.730 ;
        RECT 79.730 110.520 79.810 110.730 ;
        RECT 76.660 109.980 76.960 110.520 ;
        RECT 76.450 109.680 76.960 109.980 ;
        RECT 76.450 109.085 76.750 109.680 ;
        RECT 76.435 108.755 76.765 109.085 ;
        RECT 75.600 106.440 77.100 106.460 ;
        RECT 79.050 106.440 79.810 110.520 ;
        RECT 75.110 105.690 79.810 106.440 ;
        RECT 81.880 110.520 82.190 110.790 ;
        RECT 82.490 110.520 82.640 110.790 ;
        RECT 81.880 105.890 82.640 110.520 ;
        RECT 84.740 110.520 84.950 110.690 ;
        RECT 85.250 110.520 85.500 110.690 ;
        RECT 84.740 106.100 85.500 110.520 ;
        RECT 87.135 109.070 87.465 109.085 ;
        RECT 129.110 109.070 129.410 110.520 ;
        RECT 87.135 108.770 95.540 109.070 ;
        RECT 101.150 108.770 129.410 109.070 ;
        RECT 87.135 108.755 87.465 108.770 ;
        RECT 95.240 108.475 95.540 108.770 ;
        RECT 95.240 108.100 95.540 108.175 ;
        RECT 101.210 108.100 101.510 108.770 ;
        RECT 95.240 107.890 101.510 108.100 ;
        RECT 95.250 107.800 101.510 107.890 ;
        RECT 75.110 105.610 79.550 105.690 ;
        RECT 63.950 96.370 73.460 100.660 ;
        RECT 75.600 100.080 77.100 105.610 ;
        RECT 80.920 101.970 82.860 105.890 ;
        RECT 79.320 101.220 82.860 101.970 ;
        RECT 79.320 100.520 81.980 101.220 ;
        RECT 84.490 100.750 86.190 106.100 ;
        RECT 101.210 104.135 101.510 107.800 ;
        RECT 101.195 103.805 101.525 104.135 ;
        RECT 74.930 97.420 77.620 100.080 ;
        RECT 79.300 97.860 81.990 100.520 ;
        RECT 83.090 97.550 86.500 100.750 ;
        RECT 87.460 94.840 113.050 100.460 ;
        RECT 101.200 88.890 101.530 89.220 ;
        RECT 101.215 77.450 101.515 88.890 ;
        RECT 86.750 76.560 111.620 77.450 ;
        RECT 86.750 76.120 111.840 76.560 ;
        RECT 86.640 74.910 111.840 76.120 ;
        RECT 75.870 72.535 76.390 73.530 ;
        RECT 66.325 52.925 85.935 72.535 ;
        RECT 74.820 50.935 77.030 52.925 ;
        RECT 66.325 31.325 85.935 50.935 ;
        RECT 74.820 29.335 77.030 31.325 ;
        RECT 66.325 9.725 85.935 29.335 ;
        RECT 74.820 7.160 77.030 9.725 ;
        RECT 86.640 9.150 88.850 74.910 ;
        RECT 98.930 72.535 99.450 73.530 ;
        RECT 89.385 52.925 108.995 72.535 ;
        RECT 97.250 50.935 99.460 52.925 ;
        RECT 89.385 31.325 108.995 50.935 ;
        RECT 97.250 29.335 99.460 31.325 ;
        RECT 89.385 9.725 108.995 29.335 ;
        RECT 87.270 8.730 87.790 9.150 ;
        RECT 97.250 7.610 99.460 9.725 ;
        RECT 109.630 9.590 111.840 74.910 ;
        RECT 110.330 8.730 110.850 9.590 ;
        RECT 86.140 7.160 113.050 7.610 ;
        RECT 74.820 4.290 113.050 7.160 ;
        RECT 74.820 3.840 77.030 4.290 ;
        RECT 86.140 4.240 113.050 4.290 ;
        RECT 86.140 3.840 132.360 4.240 ;
  END
END tt_um_matt_divider_test
END LIBRARY

