VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_mingkaic1_stack_machine
  CLASS BLOCK ;
  FOREIGN tt_um_mingkaic1_stack_machine ;
  ORIGIN 0.000 0.000 ;
  SIZE 168.360 BY 225.760 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 42.670 2.480 44.270 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 83.380 2.480 84.980 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 124.090 2.480 125.690 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 164.800 2.480 166.400 223.280 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.315 2.480 23.915 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.025 2.480 64.625 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 103.735 2.480 105.335 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 144.445 2.480 146.045 223.280 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 145.670 224.760 145.970 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 148.430 224.760 148.730 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 142.910 224.760 143.210 225.760 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 137.390 224.760 137.690 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 134.630 224.760 134.930 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 131.870 224.760 132.170 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 126.350 224.760 126.650 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 123.590 224.760 123.890 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 120.830 224.760 121.130 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 115.310 224.760 115.610 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.550 224.760 112.850 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 109.790 224.760 110.090 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 104.270 224.760 104.570 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 101.510 224.760 101.810 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 98.750 224.760 99.050 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.070 224.760 49.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.310 224.760 46.610 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 43.550 224.760 43.850 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.030 224.760 38.330 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.270 224.760 35.570 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 32.510 224.760 32.810 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 71.150 224.760 71.450 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 68.390 224.760 68.690 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 65.630 224.760 65.930 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 60.110 224.760 60.410 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 57.350 224.760 57.650 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 54.590 224.760 54.890 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met4 ;
        RECT 93.230 224.760 93.530 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.462000 ;
    PORT
      LAYER met4 ;
        RECT 90.470 224.760 90.770 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met4 ;
        RECT 87.710 224.760 88.010 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met4 ;
        RECT 82.190 224.760 82.490 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.462000 ;
    PORT
      LAYER met4 ;
        RECT 79.430 224.760 79.730 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met4 ;
        RECT 76.670 224.760 76.970 225.760 ;
    END
  END uo_out[7]
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 165.600 223.125 ;
      LAYER met1 ;
        RECT 1.450 2.480 168.290 225.720 ;
      LAYER met2 ;
        RECT 1.480 2.535 168.260 225.750 ;
      LAYER met3 ;
        RECT 8.345 2.555 167.835 224.225 ;
      LAYER met4 ;
        RECT 9.495 224.360 32.110 224.760 ;
        RECT 33.210 224.360 34.870 224.760 ;
        RECT 35.970 224.360 37.630 224.760 ;
        RECT 38.730 224.360 40.390 224.760 ;
        RECT 41.490 224.360 43.150 224.760 ;
        RECT 44.250 224.360 45.910 224.760 ;
        RECT 47.010 224.360 48.670 224.760 ;
        RECT 49.770 224.360 51.430 224.760 ;
        RECT 52.530 224.360 54.190 224.760 ;
        RECT 55.290 224.360 56.950 224.760 ;
        RECT 58.050 224.360 59.710 224.760 ;
        RECT 60.810 224.360 62.470 224.760 ;
        RECT 63.570 224.360 65.230 224.760 ;
        RECT 66.330 224.360 67.990 224.760 ;
        RECT 69.090 224.360 70.750 224.760 ;
        RECT 71.850 224.360 73.510 224.760 ;
        RECT 74.610 224.360 76.270 224.760 ;
        RECT 77.370 224.360 79.030 224.760 ;
        RECT 80.130 224.360 81.790 224.760 ;
        RECT 82.890 224.360 84.550 224.760 ;
        RECT 85.650 224.360 87.310 224.760 ;
        RECT 88.410 224.360 90.070 224.760 ;
        RECT 91.170 224.360 92.830 224.760 ;
        RECT 93.930 224.360 95.590 224.760 ;
        RECT 96.690 224.360 98.350 224.760 ;
        RECT 99.450 224.360 101.110 224.760 ;
        RECT 102.210 224.360 103.870 224.760 ;
        RECT 104.970 224.360 106.630 224.760 ;
        RECT 107.730 224.360 109.390 224.760 ;
        RECT 110.490 224.360 112.150 224.760 ;
        RECT 113.250 224.360 114.910 224.760 ;
        RECT 116.010 224.360 117.670 224.760 ;
        RECT 118.770 224.360 120.430 224.760 ;
        RECT 121.530 224.360 123.190 224.760 ;
        RECT 124.290 224.360 125.950 224.760 ;
        RECT 127.050 224.360 128.710 224.760 ;
        RECT 129.810 224.360 131.470 224.760 ;
        RECT 132.570 224.360 134.230 224.760 ;
        RECT 135.330 224.360 136.990 224.760 ;
        RECT 138.090 224.360 139.750 224.760 ;
        RECT 140.850 224.360 142.510 224.760 ;
        RECT 143.610 224.360 145.270 224.760 ;
        RECT 146.370 224.360 148.030 224.760 ;
        RECT 149.130 224.360 157.945 224.760 ;
        RECT 9.495 223.680 157.945 224.360 ;
        RECT 9.495 27.375 21.915 223.680 ;
        RECT 24.315 27.375 42.270 223.680 ;
        RECT 44.670 27.375 62.625 223.680 ;
        RECT 65.025 27.375 82.980 223.680 ;
        RECT 85.380 27.375 103.335 223.680 ;
        RECT 105.735 27.375 123.690 223.680 ;
        RECT 126.090 27.375 144.045 223.680 ;
        RECT 146.445 27.375 157.945 223.680 ;
  END
END tt_um_mingkaic1_stack_machine
END LIBRARY

