VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_urish_skullfet
  CLASS BLOCK ;
  FOREIGN tt_um_urish_skullfet ;
  ORIGIN 0.000 0.000 ;
  SIZE 157.320 BY 111.520 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 10.960 21.520 12.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 20.960 21.520 22.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 30.960 21.520 32.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.960 21.520 42.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.960 21.520 52.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.960 21.520 62.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 70.960 21.520 72.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 80.960 21.520 82.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 90.960 21.520 92.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 100.960 21.520 102.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.960 21.520 112.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.960 21.520 122.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 130.960 21.520 132.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 140.960 21.520 142.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 150.960 21.520 152.560 109.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 5.960 21.520 7.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 15.960 21.520 17.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 25.960 21.520 27.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 35.960 21.520 37.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.960 21.520 47.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 55.960 21.520 57.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 65.960 21.520 67.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 75.960 21.520 77.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 85.960 21.520 87.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 95.960 21.520 97.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 105.960 21.520 107.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 115.960 21.520 117.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.960 21.520 127.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 135.960 21.520 137.560 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 145.960 21.520 147.560 109.040 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.630 110.520 134.930 111.520 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 131.870 110.520 132.170 111.520 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 129.110 110.520 129.410 111.520 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 126.350 110.520 126.650 111.520 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 123.590 110.520 123.890 111.520 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 120.830 110.520 121.130 111.520 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 110.520 118.370 111.520 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 115.310 110.520 115.610 111.520 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.550 110.520 112.850 111.520 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 109.790 110.520 110.090 111.520 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 110.520 107.330 111.520 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 104.270 110.520 104.570 111.520 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 101.510 110.520 101.810 111.520 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 98.750 110.520 99.050 111.520 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 110.520 96.290 111.520 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.230 110.520 93.530 111.520 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.470 110.520 90.770 111.520 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 87.710 110.520 88.010 111.520 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 40.790 110.520 41.090 111.520 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 38.030 110.520 38.330 111.520 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 35.270 110.520 35.570 111.520 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 32.510 110.520 32.810 111.520 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 29.750 110.520 30.050 111.520 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 26.990 110.520 27.290 111.520 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 24.230 110.520 24.530 111.520 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 62.870 110.520 63.170 111.520 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 60.110 110.520 60.410 111.520 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 57.350 110.520 57.650 111.520 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 54.590 110.520 54.890 111.520 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 51.830 110.520 52.130 111.520 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 49.070 110.520 49.370 111.520 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 46.310 110.520 46.610 111.520 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 43.550 110.520 43.850 111.520 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 84.950 110.520 85.250 111.520 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 82.190 110.520 82.490 111.520 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 79.430 110.520 79.730 111.520 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 76.670 110.520 76.970 111.520 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 73.910 110.520 74.210 111.520 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 71.150 110.520 71.450 111.520 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 68.390 110.520 68.690 111.520 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 65.630 110.520 65.930 111.520 ;
    END
  END uo_out[7]
  OBS
      LAYER nwell ;
        RECT 2.570 104.665 154.750 107.495 ;
        RECT 2.570 99.225 154.750 102.055 ;
        RECT 2.570 93.785 19.050 96.615 ;
        RECT 2.570 88.345 19.050 91.175 ;
        RECT 2.570 82.905 19.050 85.735 ;
        RECT 2.570 79.070 19.050 80.295 ;
        RECT 2.570 77.465 154.750 79.070 ;
        RECT 2.570 72.025 154.750 74.855 ;
        RECT 2.570 66.585 154.750 69.415 ;
        RECT 2.570 61.145 19.050 63.975 ;
        RECT 2.570 55.705 19.050 58.535 ;
        RECT 2.570 50.265 19.050 53.095 ;
        RECT 2.570 44.825 154.750 47.655 ;
        RECT 2.570 39.385 154.750 42.215 ;
        RECT 2.570 33.945 154.750 36.775 ;
        RECT 2.570 28.505 154.750 31.335 ;
        RECT 2.570 23.065 37.910 25.895 ;
      LAYER li1 ;
        RECT 2.760 21.675 154.560 108.885 ;
      LAYER met1 ;
        RECT 2.760 0.000 154.560 109.040 ;
      LAYER met2 ;
        RECT 5.990 0.000 152.530 110.685 ;
      LAYER met3 ;
        RECT 5.970 0.000 152.550 110.665 ;
      LAYER met4 ;
        RECT 22.170 110.120 23.830 110.665 ;
        RECT 24.930 110.120 26.590 110.665 ;
        RECT 27.690 110.120 29.350 110.665 ;
        RECT 30.450 110.120 32.110 110.665 ;
        RECT 33.210 110.120 34.870 110.665 ;
        RECT 35.970 110.120 37.630 110.665 ;
        RECT 38.730 110.120 40.390 110.665 ;
        RECT 41.490 110.120 43.150 110.665 ;
        RECT 44.250 110.120 45.910 110.665 ;
        RECT 47.010 110.120 48.670 110.665 ;
        RECT 49.770 110.120 51.430 110.665 ;
        RECT 52.530 110.120 54.190 110.665 ;
        RECT 55.290 110.120 56.950 110.665 ;
        RECT 58.050 110.120 59.710 110.665 ;
        RECT 60.810 110.120 62.470 110.665 ;
        RECT 63.570 110.120 65.230 110.665 ;
        RECT 66.330 110.120 67.990 110.665 ;
        RECT 69.090 110.120 70.750 110.665 ;
        RECT 71.850 110.120 73.510 110.665 ;
        RECT 74.610 110.120 76.270 110.665 ;
        RECT 77.370 110.120 79.030 110.665 ;
        RECT 80.130 110.120 81.790 110.665 ;
        RECT 82.890 110.120 84.550 110.665 ;
        RECT 85.650 110.120 87.310 110.665 ;
        RECT 88.410 110.120 90.070 110.665 ;
        RECT 91.170 110.120 92.830 110.665 ;
        RECT 93.930 110.120 95.590 110.665 ;
        RECT 96.690 110.120 98.350 110.665 ;
        RECT 99.450 110.120 101.110 110.665 ;
        RECT 102.210 110.120 103.870 110.665 ;
        RECT 104.970 110.120 106.630 110.665 ;
        RECT 107.730 110.120 109.390 110.665 ;
        RECT 110.490 110.120 112.150 110.665 ;
        RECT 113.250 110.120 114.910 110.665 ;
        RECT 116.010 110.120 117.670 110.665 ;
        RECT 118.770 110.120 120.430 110.665 ;
        RECT 121.530 110.120 123.190 110.665 ;
        RECT 124.290 110.120 125.950 110.665 ;
        RECT 127.050 110.120 128.710 110.665 ;
        RECT 21.455 109.440 129.425 110.120 ;
        RECT 22.960 21.120 25.560 109.440 ;
        RECT 27.960 21.120 30.560 109.440 ;
        RECT 32.960 21.120 35.560 109.440 ;
        RECT 37.960 21.120 40.560 109.440 ;
        RECT 42.960 21.120 45.560 109.440 ;
        RECT 47.960 21.120 50.560 109.440 ;
        RECT 52.960 21.120 55.560 109.440 ;
        RECT 57.960 21.120 60.560 109.440 ;
        RECT 62.960 21.120 65.560 109.440 ;
        RECT 67.960 21.120 70.560 109.440 ;
        RECT 72.960 21.120 75.560 109.440 ;
        RECT 77.960 21.120 80.560 109.440 ;
        RECT 82.960 21.120 85.560 109.440 ;
        RECT 87.960 21.120 90.560 109.440 ;
        RECT 92.960 21.120 95.560 109.440 ;
        RECT 97.960 21.120 100.560 109.440 ;
        RECT 102.960 21.120 105.560 109.440 ;
        RECT 107.960 21.120 110.560 109.440 ;
        RECT 112.960 21.120 115.560 109.440 ;
        RECT 117.960 21.120 120.560 109.440 ;
        RECT 122.960 21.120 125.560 109.440 ;
        RECT 127.960 21.120 129.425 109.440 ;
        RECT 21.455 0.000 129.425 21.120 ;
  END
END tt_um_urish_skullfet
END LIBRARY

